module rename();

endmoudle
