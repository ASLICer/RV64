module arbiter#(
    parameter OP = `R_TYPE,
    parameter OPCODE_WIDTH = 7,
    parameter REQ = 1,
    parameter AGE = 5
)(

);

endmodule